module ALU 
#
(
parameter WIDTH = 8
)
(
    input clk,
	input rstn,
    input [WIDTH-1:0] A,    // 16-bit input A
    input [WIDTH-1:0] B,    // 16-bit input B 
    input EN,
    input [3:0] ALU_FUN,
    output reg [2*WIDTH-1:0] ALU_OUT,
	output reg OUT_Valid
//    output reg Carry_Flag,
//    output reg Arith_flag, Logic_flag, CMP_flag,Shift_flag
);
//Carry_Flag = (A>B)? 1'b0:1'b1 ;
reg[2*WIDTH-1:0] D1;
reg carry_comb;
always @(posedge clk or negedge rstn) begin
	if (!rstn) begin
		ALU_OUT <= {2*WIDTH{1'b0}};
		OUT_Valid <= 1'b0;
		//Carry_Flag <= 1'b0;
	end
	else begin
	   if (EN) begin
	       ALU_OUT <= D1;
	       OUT_Valid <= 1'b1;
	       //Carry_Flag <= carry_comb;
	   end	
	   else begin
	      	ALU_OUT <= {2*WIDTH{1'b0}};
            OUT_Valid <= 1'b0;
            //Carry_Flag <= 1'b0;
	   end
	end
end
always @(*) begin
    //Carry_Flag = 0;
//	carry_comb = 0;
//    Arith_flag = 0;
//    Logic_flag = 0;
//    CMP_flag = 0;
//    Shift_flag = 0;
	D1 = 0;
    case (ALU_FUN)
        4'b0000: begin D1 = A + B; end//Arith_flag = 1; end // Addition            
        4'b0001: begin D1 = A - B; end//Arith_flag = 1; end // Subtraction
        4'b0010: begin D1 = A * B; end//Arith_flag = 1;end    // Bitwise AND
        4'b0011: begin D1 = A / B; end//Arith_flag = 1;end    // Bitwise OR
        4'b0100: begin D1 = A & B; end//Logic_flag = 1;end    // Bitwise XOR
        4'b0101: begin D1 = A | B; end//Logic_flag = 1;end
        4'b0110: begin D1 = ~(A & B); end//Logic_flag = 1;end
        4'b0111: begin D1 = ~(A | B); end//Logic_flag = 1;end
        4'b1000: begin D1 = A ^ B; end//Logic_flag = 1;end
        4'b1001: begin D1 =~(A ^ B); end//Logic_flag = 1;end
        4'b1010: begin D1 =(A==B)? 17'd1:17'd0;end //CMP_flag = 1; end 
        4'b1011: begin D1 =(A>B)? 17'd2:17'd0; end//CMP_flag = 1; end
        4'b1100: begin D1 =(A<B)? 17'd3:17'd0; end//CMP_flag = 1; end      // Bitwise NOT (only A)
        4'b1101: begin D1 = A >> 1;end //Shift_flag = 1;end   // Logical left shift
        4'b1110: begin D1 = A << 1; end//Shift_flag = 1;end   // Logical right shift
        default: begin D1 = 16'd0; end // Default case if no match
    endcase
end

    // ALU functionality to be implemented here
endmodule